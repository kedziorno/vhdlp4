library ieee;
use ieee.std_logic_1164.all;
use STD.textio.all;
use ieee.std_logic_textio.all;

package p_package is
--file file_RESULTS : text open write_mode is "output_results.txt";
end package p_package;

package body p_package is
end package body p_package;
