--
-- Definition of a single port ROM for KCPSM3 program defined by crccalc.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity crccalc is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end crccalc;
--
architecture low_level_definition of crccalc is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "1D700198AC801C70E7521730E6321620E5501510E43214004310420841044002";
attribute INIT_01 of ram_1024_x_18  : label is "1D70FCD00194AD081D70FCD00193AD101D70FCD00192AD201D70FCD00191AD40";
attribute INIT_02 of ram_1024_x_18  : label is "AD081D50FCD00190AD801D50FCD00190AD801D60FCD0AD011D70FCD00D0EAD02";
attribute INIT_03 of ram_1024_x_18  : label is "DBC001A0FCD00193AD201D40FCD00D0EAD011D50FCD00D0EAD021D50FCD00194";
attribute INIT_04 of ram_1024_x_18  : label is "1D70FCD00194AD081D70FCD00193AD101D70FCD00192AD201D700199AC401C70";
attribute INIT_05 of ram_1024_x_18  : label is "1D50FCD00191AD401D60FCD00190AD801D60FCD00D0EAD011D70FCD00195AD04";
attribute INIT_06 of ram_1024_x_18  : label is "AD101D40FCD00190AD801D40FCD0AD011D50FCD00195AD041D50FCD00191AD40";
attribute INIT_07 of ram_1024_x_18  : label is "1D70FCD00193AD101D70FCD00192AD201D700198AC801C70DBC001A1FCD00193";
attribute INIT_08 of ram_1024_x_18  : label is "1D60FCD00190AD801D60FCD00D0EAD201D70FCD00195AD401D70FCD00194AD08";
attribute INIT_09 of ram_1024_x_18  : label is "1D40FCD00D0EAD201D50FCD00192AD201D50FCD00192AD201D60FCD00191AD40";
attribute INIT_0A of ram_1024_x_18  : label is "0199AC401C70DBC001A2FCD00194AD081D40FCD00191AD401D40FCD00190AD80";
attribute INIT_0B of ram_1024_x_18  : label is "FCD00D0EAD021D70FCD00195AD041D70FCD00194AD081D70FCD00193AD201D70";
attribute INIT_0C of ram_1024_x_18  : label is "1D50FCD00192AD101D60FCD00192AD201D60FCD00191AD401D60FCD0AD011D70";
attribute INIT_0D of ram_1024_x_18  : label is "AD201D40FCD00192AD201D40FCD00191AD401D40FCD0AD011D50FCD00193AD10";
attribute INIT_0E of ram_1024_x_18  : label is "1D70FCD00195AD041D70FCD00194AD081D70019AAC401C70DBC001A3FCD00195";
attribute INIT_0F of ram_1024_x_18  : label is "AD101D60FCD00192AD201D60FCD00190AD801D60FCD0AD011D70FCD00D0EAD02";
attribute INIT_10 of ram_1024_x_18  : label is "AD201D40FCD00194AD801D40FCD00194AD081D50FCD00194AD081D60FCD00193";
attribute INIT_11 of ram_1024_x_18  : label is "1D700198AC801C70DBC001A4FCD00D0EAD021D40FCD00193AD101D40FCD00192";
attribute INIT_12 of ram_1024_x_18  : label is "AD801D60FCD0AD011D70FCD00D0EAD021D70FCD00195AD041D70FCD00193AD10";
attribute INIT_13 of ram_1024_x_18  : label is "AD041D60FCD00194AD081D60FCD00193AD101D60FCD00191AD401D60FCD00190";
attribute INIT_14 of ram_1024_x_18  : label is "AD081D40FCD00193AD101D40FCD00191AD401D40FCD00195AD041D50FCD00195";
attribute INIT_15 of ram_1024_x_18  : label is "AD101D70FCD00192AD201D700198AC801C70DBC001A5FCD0AD011D40FCD00194";
attribute INIT_16 of ram_1024_x_18  : label is "AD041D60FCD00194AD081D60FCD00192AD201D60FCD00191AD401D60FCD00193";
attribute INIT_17 of ram_1024_x_18  : label is "AD011D50FCD00194AD081D50FCD00190AD801D50FCD00D0EAD021D60FCD00195";
attribute INIT_18 of ram_1024_x_18  : label is "41A8CB10CB08CB04CB02DBC00C06FCD00195AD041D40FCD00194AD081D40FCD0";
attribute INIT_19 of ram_1024_x_18  : label is "A0000C0E0C0E0C0E0C0E0C0E0C0E0C0EA0000D0E0D0E0D0E0D0E0D0E0D0E0D0E";
attribute INIT_1A of ram_1024_x_18  : label is "00000000000000000000000000000000A0000C0E0C060C060C060C060C060C06";
attribute INIT_1B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_20 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_21 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_22 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_23 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_24 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_25 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_26 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_27 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_28 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_29 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_30 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_31 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_32 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_33 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "0C0C303303000C0C0C0C080C0C0C0C3033020203030300080C0C0C0C30000000";
attribute INITP_01 of ram_1024_x_18 : label is "030300080C0C30330303000C0C0C0C0020303030C0CC0C0C080C0C0C0C080C0C";
attribute INITP_02 of ram_1024_x_18 : label is "0303020303030303030C0C03030303030303030300080C0C3032030303030303";
attribute INITP_03 of ram_1024_x_18 : label is "00000000000000000000000000000000000000000000AAAAAAAAAAAAEA88C0C0";
attribute INITP_04 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_05 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_06 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_07 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"1D700198AC801C70E7521730E6321620E5501510E43214004310420841044002",
                INIT_01 => X"1D70FCD00194AD081D70FCD00193AD101D70FCD00192AD201D70FCD00191AD40",
                INIT_02 => X"AD081D50FCD00190AD801D50FCD00190AD801D60FCD0AD011D70FCD00D0EAD02",
                INIT_03 => X"DBC001A0FCD00193AD201D40FCD00D0EAD011D50FCD00D0EAD021D50FCD00194",
                INIT_04 => X"1D70FCD00194AD081D70FCD00193AD101D70FCD00192AD201D700199AC401C70",
                INIT_05 => X"1D50FCD00191AD401D60FCD00190AD801D60FCD00D0EAD011D70FCD00195AD04",
                INIT_06 => X"AD101D40FCD00190AD801D40FCD0AD011D50FCD00195AD041D50FCD00191AD40",
                INIT_07 => X"1D70FCD00193AD101D70FCD00192AD201D700198AC801C70DBC001A1FCD00193",
                INIT_08 => X"1D60FCD00190AD801D60FCD00D0EAD201D70FCD00195AD401D70FCD00194AD08",
                INIT_09 => X"1D40FCD00D0EAD201D50FCD00192AD201D50FCD00192AD201D60FCD00191AD40",
                INIT_0A => X"0199AC401C70DBC001A2FCD00194AD081D40FCD00191AD401D40FCD00190AD80",
                INIT_0B => X"FCD00D0EAD021D70FCD00195AD041D70FCD00194AD081D70FCD00193AD201D70",
                INIT_0C => X"1D50FCD00192AD101D60FCD00192AD201D60FCD00191AD401D60FCD0AD011D70",
                INIT_0D => X"AD201D40FCD00192AD201D40FCD00191AD401D40FCD0AD011D50FCD00193AD10",
                INIT_0E => X"1D70FCD00195AD041D70FCD00194AD081D70019AAC401C70DBC001A3FCD00195",
                INIT_0F => X"AD101D60FCD00192AD201D60FCD00190AD801D60FCD0AD011D70FCD00D0EAD02",
                INIT_10 => X"AD201D40FCD00194AD801D40FCD00194AD081D50FCD00194AD081D60FCD00193",
                INIT_11 => X"1D700198AC801C70DBC001A4FCD00D0EAD021D40FCD00193AD101D40FCD00192",
                INIT_12 => X"AD801D60FCD0AD011D70FCD00D0EAD021D70FCD00195AD041D70FCD00193AD10",
                INIT_13 => X"AD041D60FCD00194AD081D60FCD00193AD101D60FCD00191AD401D60FCD00190",
                INIT_14 => X"AD081D40FCD00193AD101D40FCD00191AD401D40FCD00195AD041D50FCD00195",
                INIT_15 => X"AD101D70FCD00192AD201D700198AC801C70DBC001A5FCD0AD011D40FCD00194",
                INIT_16 => X"AD041D60FCD00194AD081D60FCD00192AD201D60FCD00191AD401D60FCD00193",
                INIT_17 => X"AD011D50FCD00194AD081D50FCD00190AD801D50FCD00D0EAD021D60FCD00195",
                INIT_18 => X"41A8CB10CB08CB04CB02DBC00C06FCD00195AD041D40FCD00194AD081D40FCD0",
                INIT_19 => X"A0000C0E0C0E0C0E0C0E0C0E0C0E0C0EA0000D0E0D0E0D0E0D0E0D0E0D0E0D0E",
                INIT_1A => X"00000000000000000000000000000000A0000C0E0C060C060C060C060C060C06",
                INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",    
               INITP_00 => X"0C0C303303000C0C0C0C080C0C0C0C3033020203030300080C0C0C0C30000000",
               INITP_01 => X"030300080C0C30330303000C0C0C0C0020303030C0CC0C0C080C0C0C0C080C0C",
               INITP_02 => X"0303020303030303030C0C03030303030303030300080C0C3032030303030303",
               INITP_03 => X"00000000000000000000000000000000000000000000AAAAAAAAAAAAEA88C0C0",
               INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE crccalc.vhd
--
------------------------------------------------------------------------------------
