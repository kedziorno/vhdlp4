--
-- Definition of a single port ROM for KCPSM3 program defined by crccalc.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity crccalc is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end crccalc;
--
architecture low_level_definition of crccalc is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "CF010C0E0F071C70E7521730E6321620E5501510E43214004310420841044002";
attribute INIT_01 of ram_1024_x_18  : label is "FCD0541B2F00CF010D0E0F051D70FCD054142F00CF010D0E0F061D70540E2F00";
attribute INIT_02 of ram_1024_x_18  : label is "0D0E1D70FCD054292F00CF010D0E0F031D70FCD054222F00CF010D0E0F041D70";
attribute INIT_03 of ram_1024_x_18  : label is "543C2F00CF010D0E0F071D50FCD054352F00CF010D0E0F071D60FCD01D70FCD0";
attribute INIT_04 of ram_1024_x_18  : label is "0F041D40FCD00D0E1D50FCD00D0E1D50FCD054432F00CF010D0E0F031D50FCD0";
attribute INIT_05 of ram_1024_x_18  : label is "2F00CF010C0E0F061C70DBC054562F00CF010C0E0F07FCD054502F00CF010D0E";
attribute INIT_06 of ram_1024_x_18  : label is "1D70FCD0546A2F00CF010D0E0F041D70FCD054632F00CF010D0E0F051D70545D";
attribute INIT_07 of ram_1024_x_18  : label is "FCD00D0E1D70FCD054782F00CF010D0E0F021D70FCD054712F00CF010D0E0F03";
attribute INIT_08 of ram_1024_x_18  : label is "0F061D50FCD054892F00CF010D0E0F061D60FCD054822F00CF010D0E0F071D60";
attribute INIT_09 of ram_1024_x_18  : label is "0F071D40FCD01D50FCD054972F00CF010D0E0F021D50FCD054902F00CF010D0E";
attribute INIT_0A of ram_1024_x_18  : label is "2F00CF010C0E0F06FCD054A72F00CF010D0E0F041D40FCD054A02F00CF010D0E";
attribute INIT_0B of ram_1024_x_18  : label is "1D70FCD054BA2F00CF010D0E0F051D7054B42F00CF010C0E0F071C70DBC054AD";
attribute INIT_0C of ram_1024_x_18  : label is "0D0E0F021D70FCD054C82F00CF010D0E0F031D70FCD054C12F00CF010D0E0F04";
attribute INIT_0D of ram_1024_x_18  : label is "2F00CF010D0E0F071D60FCD054D62F00CF010D0E0F011D70FCD054CF2F00CF01";
attribute INIT_0E of ram_1024_x_18  : label is "FCD054EB2F00CF010D0E0F051D60FCD054E42F00CF010D0E0F061D60FCD054DD";
attribute INIT_0F of ram_1024_x_18  : label is "0F071D40FCD054F92F00CF010D0E0F011D50FCD054F22F00CF010D0E0F051D50";
attribute INIT_10 of ram_1024_x_18  : label is "CF010D0E0F031D40FCD055072F00CF010D0E0F061D40FCD055002F00CF010D0E";
attribute INIT_11 of ram_1024_x_18  : label is "1D70551B2F00CF010C0E0F061C70DBC055142F00CF010C0E0F05FCD0550E2F00";
attribute INIT_12 of ram_1024_x_18  : label is "0D0E0F021D70FCD055282F00CF010D0E0F031D70FCD055212F00CF010D0E0F04";
attribute INIT_13 of ram_1024_x_18  : label is "0D0E0F061D60FCD01D70FCD055362F00CF010D0E0F011D70FCD0552F2F00CF01";
attribute INIT_14 of ram_1024_x_18  : label is "2F00CF010D0E0F051D60FCD055462F00CF010D0E0F051D60FCD0553F2F00CF01";
attribute INIT_15 of ram_1024_x_18  : label is "2F00CF010D0E0F061D40FCD01D50FCD055542F00CF010D0E0F041D50FCD0554D";
attribute INIT_16 of ram_1024_x_18  : label is "FCD0556B2F00CF010D0E0F021D40FCD055642F00CF010D0E0F051D40FCD0555D";
attribute INIT_17 of ram_1024_x_18  : label is "000000000000000000000000CB10CB08CB04CB02DBC055712F00CF010C0E0F04";
attribute INIT_18 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_19 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_20 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_21 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_22 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_23 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_24 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_25 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_26 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_27 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_28 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_29 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_30 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_31 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_32 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_33 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "20D603580D603583580D60D602083580D603580083580D603580D60D60000000";
attribute INITP_01 of ram_1024_x_18 : label is "03580D603580D603580D603580D603580D60D603583580D6003580D603580D60";
attribute INITP_02 of ram_1024_x_18 : label is "000AA3583580D6035800D603580D6035800D603580D603583580D60D603580D6";
attribute INITP_03 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_04 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_05 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_06 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_07 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"CF010C0E0F071C70E7521730E6321620E5501510E43214004310420841044002",
                INIT_01 => X"FCD0541B2F00CF010D0E0F051D70FCD054142F00CF010D0E0F061D70540E2F00",
                INIT_02 => X"0D0E1D70FCD054292F00CF010D0E0F031D70FCD054222F00CF010D0E0F041D70",
                INIT_03 => X"543C2F00CF010D0E0F071D50FCD054352F00CF010D0E0F071D60FCD01D70FCD0",
                INIT_04 => X"0F041D40FCD00D0E1D50FCD00D0E1D50FCD054432F00CF010D0E0F031D50FCD0",
                INIT_05 => X"2F00CF010C0E0F061C70DBC054562F00CF010C0E0F07FCD054502F00CF010D0E",
                INIT_06 => X"1D70FCD0546A2F00CF010D0E0F041D70FCD054632F00CF010D0E0F051D70545D",
                INIT_07 => X"FCD00D0E1D70FCD054782F00CF010D0E0F021D70FCD054712F00CF010D0E0F03",
                INIT_08 => X"0F061D50FCD054892F00CF010D0E0F061D60FCD054822F00CF010D0E0F071D60",
                INIT_09 => X"0F071D40FCD01D50FCD054972F00CF010D0E0F021D50FCD054902F00CF010D0E",
                INIT_0A => X"2F00CF010C0E0F06FCD054A72F00CF010D0E0F041D40FCD054A02F00CF010D0E",
                INIT_0B => X"1D70FCD054BA2F00CF010D0E0F051D7054B42F00CF010C0E0F071C70DBC054AD",
                INIT_0C => X"0D0E0F021D70FCD054C82F00CF010D0E0F031D70FCD054C12F00CF010D0E0F04",
                INIT_0D => X"2F00CF010D0E0F071D60FCD054D62F00CF010D0E0F011D70FCD054CF2F00CF01",
                INIT_0E => X"FCD054EB2F00CF010D0E0F051D60FCD054E42F00CF010D0E0F061D60FCD054DD",
                INIT_0F => X"0F071D40FCD054F92F00CF010D0E0F011D50FCD054F22F00CF010D0E0F051D50",
                INIT_10 => X"CF010D0E0F031D40FCD055072F00CF010D0E0F061D40FCD055002F00CF010D0E",
                INIT_11 => X"1D70551B2F00CF010C0E0F061C70DBC055142F00CF010C0E0F05FCD0550E2F00",
                INIT_12 => X"0D0E0F021D70FCD055282F00CF010D0E0F031D70FCD055212F00CF010D0E0F04",
                INIT_13 => X"0D0E0F061D60FCD01D70FCD055362F00CF010D0E0F011D70FCD0552F2F00CF01",
                INIT_14 => X"2F00CF010D0E0F051D60FCD055462F00CF010D0E0F051D60FCD0553F2F00CF01",
                INIT_15 => X"2F00CF010D0E0F061D40FCD01D50FCD055542F00CF010D0E0F041D50FCD0554D",
                INIT_16 => X"FCD0556B2F00CF010D0E0F021D40FCD055642F00CF010D0E0F051D40FCD0555D",
                INIT_17 => X"000000000000000000000000CB10CB08CB04CB02DBC055712F00CF010C0E0F04",
                INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",    
               INITP_00 => X"20D603580D603583580D60D602083580D603580083580D603580D60D60000000",
               INITP_01 => X"03580D603580D603580D603580D603580D60D603583580D6003580D603580D60",
               INITP_02 => X"000AA3583580D6035800D603580D6035800D603580D603583580D60D603580D6",
               INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE crccalc.vhd
--
------------------------------------------------------------------------------------
