--
-- Definition of a single port ROM for KCPSM3 program defined by crccalc.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity crccalc is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end crccalc;
--
architecture low_level_definition of crccalc is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "1D7001C9AC801C70E7521730E6321620E5501510E43214004310420841044002";
attribute INIT_01 of ram_1024_x_18  : label is "1D70FCD001C5AD081D70FCD001C4AD101D70FCD001C3AD201D70FCD001C2AD40";
attribute INIT_02 of ram_1024_x_18  : label is "AD081D50FCD001C1AD801D50FCD001C1AD801D60FCD0AD011D70FCD00D0EAD02";
attribute INIT_03 of ram_1024_x_18  : label is "1C70DBC001D1FCD001C3AD201D40FCD0AD011D50FCD00D0EAD021D50FCD001C5";
attribute INIT_04 of ram_1024_x_18  : label is "AD041D70FCD001C5AD081D70FCD001C4AD101D70FCD001C3AD201D7001CAAC40";
attribute INIT_05 of ram_1024_x_18  : label is "01C2AD401D50FCD001C2AD401D60FCD001C1AD801D60FCD0AD011D70FCD001C6";
attribute INIT_06 of ram_1024_x_18  : label is "FCD001C4AD101D40FCD001C1AD801D40FCD0AD011D50FCD001C6AD041D50FCD0";
attribute INIT_07 of ram_1024_x_18  : label is "01C5AD081D70FCD001C4AD101D70FCD001C3AD201D7001C9AC801C70DBC001D2";
attribute INIT_08 of ram_1024_x_18  : label is "01C2AD401D60FCD001C1AD801D60FCD00D0EAD021D70FCD001C6AD041D70FCD0";
attribute INIT_09 of ram_1024_x_18  : label is "01C1AD801D40FCD00D0EAD021D50FCD001C3AD201D50FCD001C3AD201D60FCD0";
attribute INIT_0A of ram_1024_x_18  : label is "AD101D7001CAAC401C70DBC001D3FCD001C5AD081D40FCD001C2AD401D40FCD0";
attribute INIT_0B of ram_1024_x_18  : label is "AD011D70FCD00D0EAD021D70FCD001C6AD041D70FCD001C5AD081D70FCD001C4";
attribute INIT_0C of ram_1024_x_18  : label is "01C4AD101D50FCD001C4AD101D60FCD001C3AD201D60FCD001C2AD401D60FCD0";
attribute INIT_0D of ram_1024_x_18  : label is "FCD001C6AD041D40FCD001C3AD201D40FCD001C2AD401D40FCD0AD011D50FCD0";
attribute INIT_0E of ram_1024_x_18  : label is "0D0EAD021D70FCD001C6AD041D70FCD001C5AD081D7001CBAC401C70DBC001D4";
attribute INIT_0F of ram_1024_x_18  : label is "FCD001C4AD101D60FCD001C3AD201D60FCD001C1AD801D60FCD0AD011D70FCD0";
attribute INIT_10 of ram_1024_x_18  : label is "FCD001C3AD201D40FCD001C5AD801D40FCD001C5AD081D50FCD001C5AD081D60";
attribute INIT_11 of ram_1024_x_18  : label is "01C4AD101D7001C9AC801C70DBC001D5FCD00D0EAD021D40FCD001C4AD101D40";
attribute INIT_12 of ram_1024_x_18  : label is "FCD001C1AD801D60FCD0AD011D70FCD00D0EAD021D70FCD001C6AD041D70FCD0";
attribute INIT_13 of ram_1024_x_18  : label is "FCD001C6AD041D60FCD001C5AD081D60FCD001C4AD101D60FCD001C2AD401D60";
attribute INIT_14 of ram_1024_x_18  : label is "FCD001C5AD081D40FCD001C4AD101D40FCD001C2AD401D40FCD001C6AD041D50";
attribute INIT_15 of ram_1024_x_18  : label is "FCD001C4AD101D70FCD001C3AD201D7001C9AC801C70DBC001D6FCD0AD011D40";
attribute INIT_16 of ram_1024_x_18  : label is "FCD001C6AD041D60FCD001C5AD081D60FCD001C3AD201D60FCD001C2AD401D60";
attribute INIT_17 of ram_1024_x_18  : label is "1D40FCD0AD011D50FCD001C5AD081D50FCD001C1AD801D50FCD00D0EAD021D60";
attribute INIT_18 of ram_1024_x_18  : label is "FCD001C4AD101D7001CAAC401C70DBC00C06FCD001C6AD041D40FCD001C5AD08";
attribute INIT_19 of ram_1024_x_18  : label is "FCD001C6AD041D60FCD001C4AD101D60FCD001C3AD201D60FCD001C5AD081D70";
attribute INIT_1A of ram_1024_x_18  : label is "1D40FCD001C6AD041D50FCD001C2AD401D50FCD0AD011D60FCD00D0EAD021D60";
attribute INIT_1B of ram_1024_x_18  : label is "CB10CB08CB04CB02DBC0FCD00D0EAD021D40FCD001C6AD041D40FCD001C1AD80";
attribute INIT_1C of ram_1024_x_18  : label is "0C0E0C0E0C0E0C0E0C0E0C0E0C0EA0000D0E0D0E0D0E0D0E0D0E0D0E0D0E41D9";
attribute INIT_1D of ram_1024_x_18  : label is "0000000000000000000000000000A0000C0E0C060C060C060C060C060C06A000";
attribute INIT_1E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_1F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_20 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_21 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_22 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_23 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_24 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_25 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_26 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_27 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_28 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_29 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_30 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_31 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_32 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_33 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "C0C0C303303000C0C0C0C0030303030C0CC00203030300080C0C0C0C30000000";
attribute INITP_01 of ram_1024_x_18 : label is "3030300080C0C30330303000C0C0C0C0020303030C0CC0C0C080C0C0C0C080C0";
attribute INITP_02 of ram_1024_x_18 : label is "00303020303030303030C0C03030303030303030300080C0C303203030303030";
attribute INITP_03 of ram_1024_x_18 : label is "00000000000000000002AAAAAAAAAAABAA080C0C0C0C00203030303030C08C0C";
attribute INITP_04 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_05 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_06 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_07 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"1D7001C9AC801C70E7521730E6321620E5501510E43214004310420841044002",
                INIT_01 => X"1D70FCD001C5AD081D70FCD001C4AD101D70FCD001C3AD201D70FCD001C2AD40",
                INIT_02 => X"AD081D50FCD001C1AD801D50FCD001C1AD801D60FCD0AD011D70FCD00D0EAD02",
                INIT_03 => X"1C70DBC001D1FCD001C3AD201D40FCD0AD011D50FCD00D0EAD021D50FCD001C5",
                INIT_04 => X"AD041D70FCD001C5AD081D70FCD001C4AD101D70FCD001C3AD201D7001CAAC40",
                INIT_05 => X"01C2AD401D50FCD001C2AD401D60FCD001C1AD801D60FCD0AD011D70FCD001C6",
                INIT_06 => X"FCD001C4AD101D40FCD001C1AD801D40FCD0AD011D50FCD001C6AD041D50FCD0",
                INIT_07 => X"01C5AD081D70FCD001C4AD101D70FCD001C3AD201D7001C9AC801C70DBC001D2",
                INIT_08 => X"01C2AD401D60FCD001C1AD801D60FCD00D0EAD021D70FCD001C6AD041D70FCD0",
                INIT_09 => X"01C1AD801D40FCD00D0EAD021D50FCD001C3AD201D50FCD001C3AD201D60FCD0",
                INIT_0A => X"AD101D7001CAAC401C70DBC001D3FCD001C5AD081D40FCD001C2AD401D40FCD0",
                INIT_0B => X"AD011D70FCD00D0EAD021D70FCD001C6AD041D70FCD001C5AD081D70FCD001C4",
                INIT_0C => X"01C4AD101D50FCD001C4AD101D60FCD001C3AD201D60FCD001C2AD401D60FCD0",
                INIT_0D => X"FCD001C6AD041D40FCD001C3AD201D40FCD001C2AD401D40FCD0AD011D50FCD0",
                INIT_0E => X"0D0EAD021D70FCD001C6AD041D70FCD001C5AD081D7001CBAC401C70DBC001D4",
                INIT_0F => X"FCD001C4AD101D60FCD001C3AD201D60FCD001C1AD801D60FCD0AD011D70FCD0",
                INIT_10 => X"FCD001C3AD201D40FCD001C5AD801D40FCD001C5AD081D50FCD001C5AD081D60",
                INIT_11 => X"01C4AD101D7001C9AC801C70DBC001D5FCD00D0EAD021D40FCD001C4AD101D40",
                INIT_12 => X"FCD001C1AD801D60FCD0AD011D70FCD00D0EAD021D70FCD001C6AD041D70FCD0",
                INIT_13 => X"FCD001C6AD041D60FCD001C5AD081D60FCD001C4AD101D60FCD001C2AD401D60",
                INIT_14 => X"FCD001C5AD081D40FCD001C4AD101D40FCD001C2AD401D40FCD001C6AD041D50",
                INIT_15 => X"FCD001C4AD101D70FCD001C3AD201D7001C9AC801C70DBC001D6FCD0AD011D40",
                INIT_16 => X"FCD001C6AD041D60FCD001C5AD081D60FCD001C3AD201D60FCD001C2AD401D60",
                INIT_17 => X"1D40FCD0AD011D50FCD001C5AD081D50FCD001C1AD801D50FCD00D0EAD021D60",
                INIT_18 => X"FCD001C4AD101D7001CAAC401C70DBC00C06FCD001C6AD041D40FCD001C5AD08",
                INIT_19 => X"FCD001C6AD041D60FCD001C4AD101D60FCD001C3AD201D60FCD001C5AD081D70",
                INIT_1A => X"1D40FCD001C6AD041D50FCD001C2AD401D50FCD0AD011D60FCD00D0EAD021D60",
                INIT_1B => X"CB10CB08CB04CB02DBC0FCD00D0EAD021D40FCD001C6AD041D40FCD001C1AD80",
                INIT_1C => X"0C0E0C0E0C0E0C0E0C0E0C0E0C0EA0000D0E0D0E0D0E0D0E0D0E0D0E0D0E41D9",
                INIT_1D => X"0000000000000000000000000000A0000C0E0C060C060C060C060C060C06A000",
                INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",    
               INITP_00 => X"C0C0C303303000C0C0C0C0030303030C0CC00203030300080C0C0C0C30000000",
               INITP_01 => X"3030300080C0C30330303000C0C0C0C0020303030C0CC0C0C080C0C0C0C080C0",
               INITP_02 => X"00303020303030303030C0C03030303030303030300080C0C303203030303030",
               INITP_03 => X"00000000000000000002AAAAAAAAAAABAA080C0C0C0C00203030303030C08C0C",
               INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE crccalc.vhd
--
------------------------------------------------------------------------------------
